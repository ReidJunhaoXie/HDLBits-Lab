`timescale 1ns/1ps 
module simple_wire_02( input in, output out );
   assign out = in ; 
endmodule
