`timescale 1ns/1ps

module rtl_7458_chip_07(
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );
    
    assign p1y = (p1a&p1b&p1c)|(p1d&p1e&p1f) ;
    assign p2y = (p2a&p2b)|(p2c&p2d) ;
    
endmodule