`timescale 1ns/1ps 
module not_gate_04(
    input in,
    output out
) ;
    assign out = ~in ;
endmodule