module wire_01( output out );
    assign out = 1'b1 ;
endmodule